module not_gate_dt (
	input a,
	output y
);
	assign y = ~a;
endmodule